-- BMP format V4HEADER